`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/03/25 15:59:18
// Design Name: 
// Module Name: test_tcam
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test();

reg clk;
reg reset;
reg [2047:0] message;



initial
begin
clk=0;
forever 
#5 clk=!clk;
end

initial
begin
reset=1;
#10 reset=0;
#10 reset=1;
end

top u_top(
.message(message),
.clk(clk),
.reset(reset)
);    

initial begin



message=2048'h7a7ac0a8c8010000000000338100000081000000884700064140450000400001000040016948c0a8c821c0a8c70108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#30
message=2048'h7a7ac0a8c801000000000033810000000800450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h01005e000009000000000033080046000024000100000111a544c0a8c821e0000009fdafad0002080208000c91f0010200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
/*
message=2048'h7a7ac0a8c80100000000003386dd6000000000340040fe800000000000000000000000000033fe8000000000000000000000000000013c000000000000002b000000000000002c000000000000000600000000000000000700070000000000000000500227108b8f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#30
message=2048'h7a7ac0a8c80100000000003386dd6000000000383c40fe800000000000000000000000000034fe8000000000000000000000000000022b020101140000010e2544142431231211212221212121002c000000000000003c000000000000001100000000000000020802080008fe980000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h01005e000009000000000033080046000024000100000111a544c0a8c821e0000009fdafad0002080208000c91f0010200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c801000000000033884700000040000000400000004000000140450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c8010000000000338100000081000000884700000040000000400000004000000140450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003381000000810000000800450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c8010000000000330800450000400001000240016946c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c8010000000000330800450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c801000000000033080600010800060400010000000000aac0a8c821000000000000c0a8c80100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003381000000080600010800060400010000000000aac0441421000000000000bf5c1401000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c8010000000000338100000081000000080600010800060400010000000000aa0c0802210000000000005b0200010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003308004500001c000100004011695cc0a8c821c0a8c801020802080008ea5900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;



message=2048'h7a7ac0a8c80100000000003386dd6000000000200040fe800000000000000000000000000033fe8000000000000000000000000000011102010ff0dfa0fa00f0df00000000000000000000000000020802080008fe980000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#30

message=2048'h7a7ac0a8c80100000000003386dd60000000002c0040fe800000000000000000000000000033fe8000000000000000000000000000010602010ff0dfa0fa00f0df00000000000000000000000000000700070000000000000000500227108b8f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003386dd6000000000140640fe800000000000000000000000000033fe800000000000000000000000000001000700070000000000000000500227108b8f000000000000000700070000000000000000500227108b8f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003308004b000040000100004006aa4ec0a8c821c0a8c801a0df00f0a0dfda00f00000f0d0a0fa0000b0f0000000f000000700070000000000000000500227107750000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c801000000000033080045000028000100004006695bc0a8c821c0a8c80100070007000000000000000050022710775000000000f000000700070000000000000000500227107750000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003308004500004a000100004032690dc0a8c821c0a8c801123456780000000008005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003308004a00005e000100004032e78cc0a8c821c0a8c801d0a0fa00000000f0af00000000fb00df00000000123456780000000008005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003386dd6000000000363240fe800000000000000000000000000033fe800000000000000000000000000001123456780000000008005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003386dd60000000003e0040fe800000000000000000000000000033fe8000000000000000000000000000013200000000000000123456780000000008005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
message=2048'h7a7ac0a8c80100000000003381000000810000000800450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#30
message=2048'h7a7ac0a8c801000000000033884700064140450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c801000000000033080045000028000100004006695bc0a8c821c0a8c801000700070000000000000000500227107750000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c80100000000003386dd6000000000363240fe800000000000000000000000000033fe800000000000000000000000000001000000010000000008005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c801000000000033810000000800450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#10
message=2048'h7a7ac0a8c801000000000033884700000040000000400000004000000140450000400001000040016948c0a8c821c0a8c80108005f5d00010001313233343536373839306162636465666768696a6b6c6d6e6f707172737475767778797a000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
*/
end
    

endmodule